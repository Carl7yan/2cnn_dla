`ifndef TESTBENCH_PKG__SV
`define TESTBENCH_PKG__SV

package testbench_pkg;
    import uvm_pkg::*;
    import PKG_dla_typedef::*;
    `include "driver_cbs.sv"
    `include "driver_cbs_coverage.sv"
    `include "transaction.sv"

    `include "kpe_driver.sv"
    `include "kpe_mon.sv"
    `include "kpe_sequencer.sv"
    `include "in_agt.sv"
    `include "out_agt.sv"

    `include "kpe_model.sv"
    `include "kpe_scoreboard.sv"
    `include "kpe_env.sv"
    `include "virtual_sequencer.sv"
    `include "base_test.sv"
    `include "case0_sequence.sv"
    `include "case1_sequence.sv"
    `include "case2_sequence.sv"
    `include "case3_sequence.sv"
    `include "case4_sequence.sv"
    `include "my_case.sv"

endpackage
`endif
