`ifndef REG_MODEL_PKG__SV
`define REG_MODEL_PKG__SV

package reg_model_pkg;
    import uvm_pkg::*;
    import reg_field_pkg::*;
    import reg_block_pkg::*;
    `include "reg_model.sv"
endpackage
`endif 